library ieee;
use ieee.std_logic_1164.all;

entity TFF is
port( din: in std_logic;
clk: in std_logic;
rst: in std_logic;
dout: out std_logic);
end TFF;

architecture behavioral of TFF is
begin
process(rst,clk,din)
begin
if (rst='1') then
dout<='0';
elsif(rising_edge(clk)) then
dout<=not din;
end if;
end process;

end behavioral;
